VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SRAM_32x1024_2P
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 278.464 BY 66.880 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.568 0.000 263.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 263.568 0.000 263.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 263.568 0.000 263.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 263.568 0.000 263.720 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.016 0.000 252.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 252.016 0.000 252.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 252.016 0.000 252.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 252.016 0.000 252.168 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.464 0.000 240.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 240.464 0.000 240.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 240.464 0.000 240.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 240.464 0.000 240.616 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.912 0.000 229.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 228.912 0.000 229.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 228.912 0.000 229.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 228.912 0.000 229.064 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.608 0.000 228.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 228.608 0.000 228.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 228.608 0.000 228.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 228.608 0.000 228.760 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.304 0.000 228.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 228.304 0.000 228.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 228.304 0.000 228.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 228.304 0.000 228.456 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.000 0.000 228.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 228.000 0.000 228.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 228.000 0.000 228.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 228.000 0.000 228.152 0.152 ;
    END
  END O1[0]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.448 0.000 216.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 216.448 0.000 216.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 216.448 0.000 216.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 216.448 0.000 216.600 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.984 0.000 204.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 203.984 0.000 204.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 203.984 0.000 204.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 203.984 0.000 204.136 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.680 0.000 203.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 203.680 0.000 203.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 203.680 0.000 203.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 203.680 0.000 203.832 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.376 0.000 203.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 203.376 0.000 203.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 203.376 0.000 203.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 203.376 0.000 203.528 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.072 0.000 203.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 203.072 0.000 203.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 203.072 0.000 203.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 203.072 0.000 203.224 0.152 ;
    END
  END O1[8]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.520 0.000 191.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 191.520 0.000 191.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 191.520 0.000 191.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 191.520 0.000 191.672 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.216 0.000 191.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 191.216 0.000 191.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 191.216 0.000 191.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 191.216 0.000 191.368 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.912 0.000 191.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.912 0.000 191.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.912 0.000 191.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.912 0.000 191.064 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
  END O1[12]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.056 0.000 179.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 179.056 0.000 179.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 179.056 0.000 179.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.056 0.000 179.208 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.752 0.000 178.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 178.752 0.000 178.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 178.752 0.000 178.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 178.752 0.000 178.904 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.448 0.000 178.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 178.448 0.000 178.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 178.448 0.000 178.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 178.448 0.000 178.600 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.144 0.000 178.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 178.144 0.000 178.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 178.144 0.000 178.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 178.144 0.000 178.296 0.152 ;
    END
  END O1[16]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.592 0.000 166.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 166.592 0.000 166.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 166.592 0.000 166.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 166.592 0.000 166.744 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.288 0.000 166.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 166.288 0.000 166.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 166.288 0.000 166.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 166.288 0.000 166.440 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.984 0.000 166.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 165.984 0.000 166.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 165.984 0.000 166.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 165.984 0.000 166.136 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.680 0.000 165.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 165.680 0.000 165.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 165.680 0.000 165.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 165.680 0.000 165.832 0.152 ;
    END
  END O1[20]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
  END O1[24]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.752 0.000 140.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 140.752 0.000 140.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 140.752 0.000 140.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.752 0.000 140.904 0.152 ;
    END
  END O1[28]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 58.520 278.464 58.672 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 58.520 278.464 58.672 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 58.520 278.464 58.672 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 58.520 278.464 58.672 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 54.872 278.464 55.024 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 54.872 278.464 55.024 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 54.872 278.464 55.024 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 54.872 278.464 55.024 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 51.224 278.464 51.376 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 51.224 278.464 51.376 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 51.224 278.464 51.376 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 51.224 278.464 51.376 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 47.576 278.464 47.728 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 47.576 278.464 47.728 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 47.576 278.464 47.728 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 47.576 278.464 47.728 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 43.928 278.464 44.080 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 43.928 278.464 44.080 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 43.928 278.464 44.080 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 43.928 278.464 44.080 ;
    END
  END A1[4]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 40.280 278.464 40.432 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 40.280 278.464 40.432 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 40.280 278.464 40.432 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 40.280 278.464 40.432 ;
    END
  END A1[5]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 36.632 278.464 36.784 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 36.632 278.464 36.784 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 36.632 278.464 36.784 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 36.632 278.464 36.784 ;
    END
  END A1[6]

  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 32.984 278.464 33.136 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 32.984 278.464 33.136 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 32.984 278.464 33.136 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 32.984 278.464 33.136 ;
    END
  END A1[7]

  PIN A1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 29.336 278.464 29.488 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 29.336 278.464 29.488 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 29.336 278.464 29.488 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 29.336 278.464 29.488 ;
    END
  END A1[8]

  PIN A1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 25.688 278.464 25.840 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 25.688 278.464 25.840 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 25.688 278.464 25.840 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 25.688 278.464 25.840 ;
    END
  END A1[9]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.896 0.000 15.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.896 0.000 15.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.896 0.000 15.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.896 0.000 15.048 0.152 ;
    END
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.448 0.000 26.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.448 0.000 26.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.448 0.000 26.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.448 0.000 26.600 0.152 ;
    END
  END CSB2

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
  END I2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
  END I2[1]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
  END I2[2]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
  END I2[3]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
  END I2[4]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
  END I2[5]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
  END I2[6]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
  END I2[7]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.928 0.000 63.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.928 0.000 63.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.928 0.000 63.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.928 0.000 63.080 0.152 ;
    END
  END I2[8]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
  END I2[9]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
  END I2[10]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
  END I2[11]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
  END I2[12]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
  END I2[13]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
  END I2[14]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
  END I2[15]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
  END I2[16]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
  END I2[17]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
  END I2[18]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
  END I2[19]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
  END I2[20]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
  END I2[21]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
  END I2[22]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
  END I2[23]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
  END I2[24]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.088 0.000 113.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.088 0.000 113.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.088 0.000 113.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.088 0.000 113.240 0.152 ;
    END
  END I2[25]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.392 0.000 113.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.392 0.000 113.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.392 0.000 113.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.392 0.000 113.544 0.152 ;
    END
  END I2[26]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.696 0.000 113.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.696 0.000 113.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.696 0.000 113.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.696 0.000 113.848 0.152 ;
    END
  END I2[27]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
  END I2[28]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
  END I2[29]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
  END I2[30]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
  END I2[31]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 58.520 0.152 58.672 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 58.520 0.152 58.672 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 58.520 0.152 58.672 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 58.520 0.152 58.672 ;
    END
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 54.872 0.152 55.024 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 54.872 0.152 55.024 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 54.872 0.152 55.024 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 54.872 0.152 55.024 ;
    END
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 51.224 0.152 51.376 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 51.224 0.152 51.376 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 51.224 0.152 51.376 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 51.224 0.152 51.376 ;
    END
  END A2[2]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 47.576 0.152 47.728 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 47.576 0.152 47.728 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 47.576 0.152 47.728 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 47.576 0.152 47.728 ;
    END
  END A2[3]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 43.928 0.152 44.080 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 43.928 0.152 44.080 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 43.928 0.152 44.080 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 43.928 0.152 44.080 ;
    END
  END A2[4]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 40.280 0.152 40.432 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 40.280 0.152 40.432 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 40.280 0.152 40.432 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 40.280 0.152 40.432 ;
    END
  END A2[5]

  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 36.632 0.152 36.784 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 36.632 0.152 36.784 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 36.632 0.152 36.784 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 36.632 0.152 36.784 ;
    END
  END A2[6]

  PIN A2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 32.984 0.152 33.136 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 32.984 0.152 33.136 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 32.984 0.152 33.136 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 32.984 0.152 33.136 ;
    END
  END A2[7]

  PIN A2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 29.336 0.152 29.488 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 29.336 0.152 29.488 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 29.336 0.152 29.488 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 29.336 0.152 29.488 ;
    END
  END A2[8]

  PIN A2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 25.688 0.152 25.840 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 25.688 0.152 25.840 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 25.688 0.152 25.840 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 25.688 0.152 25.840 ;
    END
  END A2[9]

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 16.720 0.152 16.872 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 16.720 0.152 16.872 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 16.720 0.152 16.872 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 16.720 0.152 16.872 ;
    END
  END WEB2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 64.880 7.195 66.880 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 64.880 7.195 66.880 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 64.880 7.195 66.880 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 64.880 9.915 66.880 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 64.880 9.915 66.880 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 64.880 9.915 66.880 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 263.872 0.000 278.464 0.304 ;
      RECT 252.320 0.000 263.416 0.304 ;
      RECT 240.768 0.000 251.864 0.304 ;
      RECT 229.216 0.000 240.312 0.304 ;
      RECT 216.752 0.000 227.848 0.304 ;
      RECT 204.288 0.000 215.384 0.304 ;
      RECT 191.824 0.000 202.920 0.304 ;
      RECT 179.360 0.000 190.456 0.304 ;
      RECT 166.896 0.000 177.992 0.304 ;
      RECT 154.432 0.000 165.528 0.304 ;
      RECT 141.968 0.000 153.064 0.304 ;
      RECT 278.160 58.824 278.464 64.728 ;
      RECT 278.160 55.176 278.464 58.368 ;
      RECT 278.160 51.528 278.464 54.720 ;
      RECT 278.160 47.880 278.464 51.072 ;
      RECT 278.160 44.232 278.464 47.424 ;
      RECT 278.160 40.584 278.464 43.776 ;
      RECT 278.160 36.936 278.464 40.128 ;
      RECT 278.160 33.288 278.464 36.480 ;
      RECT 278.160 29.640 278.464 32.832 ;
      RECT 278.160 25.992 278.464 29.184 ;
      RECT 278.160 17.024 278.464 25.536 ;
      RECT 278.160 0.304 278.464 16.568 ;
      RECT 0.000 0.000 14.744 0.304 ;
      RECT 15.200 0.000 26.296 0.304 ;
      RECT 26.752 0.000 37.848 0.304 ;
      RECT 39.216 0.000 50.312 0.304 ;
      RECT 51.680 0.000 62.776 0.304 ;
      RECT 64.144 0.000 75.240 0.304 ;
      RECT 76.608 0.000 87.704 0.304 ;
      RECT 89.072 0.000 100.168 0.304 ;
      RECT 101.536 0.000 112.632 0.304 ;
      RECT 114.000 0.000 125.096 0.304 ;
      RECT 126.464 0.000 140.600 0.304 ;
      RECT 0.000 58.824 0.304 64.728 ;
      RECT 0.000 55.176 0.304 58.368 ;
      RECT 0.000 51.528 0.304 54.720 ;
      RECT 0.000 47.880 0.304 51.072 ;
      RECT 0.000 44.232 0.304 47.424 ;
      RECT 0.000 40.584 0.304 43.776 ;
      RECT 0.000 36.936 0.304 40.128 ;
      RECT 0.000 33.288 0.304 36.480 ;
      RECT 0.000 29.640 0.304 32.832 ;
      RECT 0.000 25.992 0.304 29.184 ;
      RECT 0.000 17.024 0.304 25.536 ;
      RECT 0.000 0.304 0.304 16.568 ;
      RECT 0.000 64.728 5.043 66.880 ;
      RECT 7.355 64.728 7.763 66.880 ;
      RECT 10.067 64.728 278.464 66.880 ;
      RECT 0.304 0.304 278.160 64.728 ;
    LAYER M3 ;
      RECT 263.872 0.000 278.464 0.304 ;
      RECT 252.320 0.000 263.416 0.304 ;
      RECT 240.768 0.000 251.864 0.304 ;
      RECT 229.216 0.000 240.312 0.304 ;
      RECT 216.752 0.000 227.848 0.304 ;
      RECT 204.288 0.000 215.384 0.304 ;
      RECT 191.824 0.000 202.920 0.304 ;
      RECT 179.360 0.000 190.456 0.304 ;
      RECT 166.896 0.000 177.992 0.304 ;
      RECT 154.432 0.000 165.528 0.304 ;
      RECT 141.968 0.000 153.064 0.304 ;
      RECT 278.160 58.824 278.464 64.728 ;
      RECT 278.160 55.176 278.464 58.368 ;
      RECT 278.160 51.528 278.464 54.720 ;
      RECT 278.160 47.880 278.464 51.072 ;
      RECT 278.160 44.232 278.464 47.424 ;
      RECT 278.160 40.584 278.464 43.776 ;
      RECT 278.160 36.936 278.464 40.128 ;
      RECT 278.160 33.288 278.464 36.480 ;
      RECT 278.160 29.640 278.464 32.832 ;
      RECT 278.160 25.992 278.464 29.184 ;
      RECT 278.160 17.024 278.464 25.536 ;
      RECT 278.160 0.304 278.464 16.568 ;
      RECT 0.000 0.000 14.744 0.304 ;
      RECT 15.200 0.000 26.296 0.304 ;
      RECT 26.752 0.000 37.848 0.304 ;
      RECT 39.216 0.000 50.312 0.304 ;
      RECT 51.680 0.000 62.776 0.304 ;
      RECT 64.144 0.000 75.240 0.304 ;
      RECT 76.608 0.000 87.704 0.304 ;
      RECT 89.072 0.000 100.168 0.304 ;
      RECT 101.536 0.000 112.632 0.304 ;
      RECT 114.000 0.000 125.096 0.304 ;
      RECT 126.464 0.000 140.600 0.304 ;
      RECT 0.000 58.824 0.304 64.728 ;
      RECT 0.000 55.176 0.304 58.368 ;
      RECT 0.000 51.528 0.304 54.720 ;
      RECT 0.000 47.880 0.304 51.072 ;
      RECT 0.000 44.232 0.304 47.424 ;
      RECT 0.000 40.584 0.304 43.776 ;
      RECT 0.000 36.936 0.304 40.128 ;
      RECT 0.000 33.288 0.304 36.480 ;
      RECT 0.000 29.640 0.304 32.832 ;
      RECT 0.000 25.992 0.304 29.184 ;
      RECT 0.000 17.024 0.304 25.536 ;
      RECT 0.000 0.304 0.304 16.568 ;
      RECT 0.000 64.728 5.043 66.880 ;
      RECT 7.355 64.728 7.763 66.880 ;
      RECT 10.067 64.728 278.464 66.880 ;
      RECT 0.304 0.304 278.160 64.728 ;
    LAYER M4 ;
      RECT 263.872 0.000 278.464 0.304 ;
      RECT 252.320 0.000 263.416 0.304 ;
      RECT 240.768 0.000 251.864 0.304 ;
      RECT 229.216 0.000 240.312 0.304 ;
      RECT 216.752 0.000 227.848 0.304 ;
      RECT 204.288 0.000 215.384 0.304 ;
      RECT 191.824 0.000 202.920 0.304 ;
      RECT 179.360 0.000 190.456 0.304 ;
      RECT 166.896 0.000 177.992 0.304 ;
      RECT 154.432 0.000 165.528 0.304 ;
      RECT 141.968 0.000 153.064 0.304 ;
      RECT 278.160 58.824 278.464 64.728 ;
      RECT 278.160 55.176 278.464 58.368 ;
      RECT 278.160 51.528 278.464 54.720 ;
      RECT 278.160 47.880 278.464 51.072 ;
      RECT 278.160 44.232 278.464 47.424 ;
      RECT 278.160 40.584 278.464 43.776 ;
      RECT 278.160 36.936 278.464 40.128 ;
      RECT 278.160 33.288 278.464 36.480 ;
      RECT 278.160 29.640 278.464 32.832 ;
      RECT 278.160 25.992 278.464 29.184 ;
      RECT 278.160 17.024 278.464 25.536 ;
      RECT 278.160 0.304 278.464 16.568 ;
      RECT 0.000 0.000 14.744 0.304 ;
      RECT 15.200 0.000 26.296 0.304 ;
      RECT 26.752 0.000 37.848 0.304 ;
      RECT 39.216 0.000 50.312 0.304 ;
      RECT 51.680 0.000 62.776 0.304 ;
      RECT 64.144 0.000 75.240 0.304 ;
      RECT 76.608 0.000 87.704 0.304 ;
      RECT 89.072 0.000 100.168 0.304 ;
      RECT 101.536 0.000 112.632 0.304 ;
      RECT 114.000 0.000 125.096 0.304 ;
      RECT 126.464 0.000 140.600 0.304 ;
      RECT 0.000 58.824 0.304 64.728 ;
      RECT 0.000 55.176 0.304 58.368 ;
      RECT 0.000 51.528 0.304 54.720 ;
      RECT 0.000 47.880 0.304 51.072 ;
      RECT 0.000 44.232 0.304 47.424 ;
      RECT 0.000 40.584 0.304 43.776 ;
      RECT 0.000 36.936 0.304 40.128 ;
      RECT 0.000 33.288 0.304 36.480 ;
      RECT 0.000 29.640 0.304 32.832 ;
      RECT 0.000 25.992 0.304 29.184 ;
      RECT 0.000 17.024 0.304 25.536 ;
      RECT 0.000 0.304 0.304 16.568 ;
      RECT 0.000 64.728 5.043 66.880 ;
      RECT 7.355 64.728 7.763 66.880 ;
      RECT 10.067 64.728 278.464 66.880 ;
      RECT 0.304 0.304 278.160 64.728 ;
    LAYER M5 ;
      RECT 263.872 0.000 278.464 0.304 ;
      RECT 252.320 0.000 263.416 0.304 ;
      RECT 240.768 0.000 251.864 0.304 ;
      RECT 229.216 0.000 240.312 0.304 ;
      RECT 216.752 0.000 227.848 0.304 ;
      RECT 204.288 0.000 215.384 0.304 ;
      RECT 191.824 0.000 202.920 0.304 ;
      RECT 179.360 0.000 190.456 0.304 ;
      RECT 166.896 0.000 177.992 0.304 ;
      RECT 154.432 0.000 165.528 0.304 ;
      RECT 141.968 0.000 153.064 0.304 ;
      RECT 278.160 58.824 278.464 64.728 ;
      RECT 278.160 55.176 278.464 58.368 ;
      RECT 278.160 51.528 278.464 54.720 ;
      RECT 278.160 47.880 278.464 51.072 ;
      RECT 278.160 44.232 278.464 47.424 ;
      RECT 278.160 40.584 278.464 43.776 ;
      RECT 278.160 36.936 278.464 40.128 ;
      RECT 278.160 33.288 278.464 36.480 ;
      RECT 278.160 29.640 278.464 32.832 ;
      RECT 278.160 25.992 278.464 29.184 ;
      RECT 278.160 17.024 278.464 25.536 ;
      RECT 278.160 0.304 278.464 16.568 ;
      RECT 0.000 0.000 14.744 0.304 ;
      RECT 15.200 0.000 26.296 0.304 ;
      RECT 26.752 0.000 37.848 0.304 ;
      RECT 39.216 0.000 50.312 0.304 ;
      RECT 51.680 0.000 62.776 0.304 ;
      RECT 64.144 0.000 75.240 0.304 ;
      RECT 76.608 0.000 87.704 0.304 ;
      RECT 89.072 0.000 100.168 0.304 ;
      RECT 101.536 0.000 112.632 0.304 ;
      RECT 114.000 0.000 125.096 0.304 ;
      RECT 126.464 0.000 140.600 0.304 ;
      RECT 0.000 58.824 0.304 64.728 ;
      RECT 0.000 55.176 0.304 58.368 ;
      RECT 0.000 51.528 0.304 54.720 ;
      RECT 0.000 47.880 0.304 51.072 ;
      RECT 0.000 44.232 0.304 47.424 ;
      RECT 0.000 40.584 0.304 43.776 ;
      RECT 0.000 36.936 0.304 40.128 ;
      RECT 0.000 33.288 0.304 36.480 ;
      RECT 0.000 29.640 0.304 32.832 ;
      RECT 0.000 25.992 0.304 29.184 ;
      RECT 0.000 17.024 0.304 25.536 ;
      RECT 0.000 0.304 0.304 16.568 ;
      RECT 0.000 64.728 5.043 66.880 ;
      RECT 7.355 64.728 7.763 66.880 ;
      RECT 10.067 64.728 278.464 66.880 ;
      RECT 0.304 0.304 278.160 64.728 ;
  END

END SRAM_32x1024_2P

END LIBRARY
